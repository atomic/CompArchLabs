`timescale 1ns / 1ps

module regfile(
	input clk,
	input regwrite,
	input [4:0] rr1, rr2, wr,
	input [31:0] wdata,
	output [31:0] rdata1, rdata2
);
	
	

endmodule